package soc_module_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "wb_x_uart_ref_model.sv"
	`include "wb_interconnect_ref_model.sv"
	`include "soc_scoreboard.sv"
	`include "soc_module.sv"
endpackage

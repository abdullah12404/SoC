`define UART_BASE_ADDRESS 32'h20000000
`define UART_END_ADDRESS 32'h200000FF

`define GPIO_BASE_ADDRESS 32'h20000100
`define GPIO_END_ADDRESS 32'h200001FF

`define SPI1_BASE_ADDRESS 32'h20000200
`define SPI1_END_ADDRESS 32'h2000027F

`define SPI2_BASE_ADDRESS 32'h20000280
`define SPI2_END_ADDRESS 32'h200002FF

`define I2C_BASE_ADDRESS 32'h20000300
`define I2C_END_ADDRESS 32'h200003FF


`define PTC_BASE_ADDRESS 32'h20000400
`define PTC_END_ADDRESS 32'h200004FF

`define CLINT_BASE_ADDRESS 32'h20000C00
`define CLINT_END_ADDRESS 32'h20000C0F

`define UART_BASE_ADDRESS 32'h20000000
